`timescale 1ps/1ps

module _____00003aT0( ); 
   reg clk;
   reg rst;
   reg req;
   reg ackA;
   reg ackB;
   reg ack;
   reg fill;
   wire [7:0] _00003a14;
   reg _00003a12;
   reg [0:0] _00003a13;
   wire [7:0] _00003a43;
   reg _00003a41;
   reg [0:0] _00003a42;
   wire [7:0] _00003a72;
   reg _00003a70;
   reg [0:0] _00003a71;
   reg [7:0] _00003a89;
   reg [7:0] _00003a90;
   wire [7:0] _00003a120;
   wire [7:0] _00003a121;
   reg [7:0] _00003a150;
   reg [7:0] _00003a151;
   reg [7:0] _00003a181;
   reg [7:0] _00003a182;
   reg [7:0] z0__val;
   reg [7:0] z1__val;
   wire [7:0] a0__val;
   wire [7:0] a1__val;
   reg _00003a16;
   reg [0:0] _00003a17;
   reg [7:0] _00003a18;
   reg _00003a45;
   reg [0:0] _00003a46;
   reg [7:0] _00003a47;
   reg _00003a74;
   reg [0:0] _00003a75;
   reg [7:0] _00003a76;
   reg [7:0] _00003a135;
   reg [7:0] _00003a136;
   reg [0:0] _00003a137;
   reg [7:0] val;
   wire _00003a331_00003a_00003atrig__r;
   wire _00003a331_00003a_00003atrig__w;
   reg [7:0] _00003a331_00003a_00003adbus__r;
   wire [7:0] _00003a331_00003a_00003adbus__w;
   wire [0:0] _00003a331_00003a_00003aabus__r;
   wire [0:0] _00003a331_00003a_00003aabus__w;
   reg [7:0] _00003a331_00003a_00003amem  [0:1];
   wire _00003a332_00003a_00003atrig__r;
   wire _00003a332_00003a_00003atrig__w;
   reg [7:0] _00003a332_00003a_00003adbus__r;
   wire [7:0] _00003a332_00003a_00003adbus__w;
   wire [0:0] _00003a332_00003a_00003aabus__r;
   wire [0:0] _00003a332_00003a_00003aabus__w;
   reg [7:0] _00003a332_00003a_00003amem  [0:1];
   wire _00003a333_00003a_00003atrig__r;
   wire _00003a333_00003a_00003atrig__w;
   reg [7:0] _00003a333_00003a_00003adbus__r;
   wire [7:0] _00003a333_00003a_00003adbus__w;
   wire [0:0] _00003a333_00003a_00003aabus__r;
   wire [0:0] _00003a333_00003a_00003aabus__w;
   reg [7:0] _00003a333_00003a_00003amem  [0:1];
   wire [7:0] _00003a334_00003a_00003areg__0;
   wire [7:0] _00003a334_00003a_00003areg__1;
   wire [0:0] _00003a334_00003a_00003a_00003a237_00003a_00003aabus__r;
   wire [0:0] _00003a334_00003a_00003a_00003a238_00003a_00003aabus__w;
   wire [0:0] _00003a334_00003a_00003a_00003a239_00003a_00003aabus__r;
   wire [0:0] _00003a334_00003a_00003a_00003a240_00003a_00003aabus__w;
   reg [7:0] _00003a335_00003a_00003alv0;
   reg [7:0] _00003a335_00003a_00003alv1;
   reg [7:0] _00003a335_00003a_00003aav0;
   reg [7:0] _00003a335_00003a_00003aav1;
   reg [7:0] _00003a335_00003a_00003arv;
   reg _00003a335_00003a_00003alvok0;
   reg _00003a335_00003a_00003alvok1;
   reg _00003a335_00003a_00003arvok;
   reg _00003a335_00003a_00003arun;
   wire [7:0] _00003a336_00003a_00003areg__0;
   wire [7:0] _00003a336_00003a_00003areg__1;
   wire [0:0] _00003a336_00003a_00003a_00003a268_00003a_00003aabus__r;
   wire [0:0] _00003a336_00003a_00003a_00003a269_00003a_00003aabus__w;
   wire [0:0] _00003a336_00003a_00003a_00003a270_00003a_00003aabus__r;
   wire [0:0] _00003a336_00003a_00003a_00003a271_00003a_00003aabus__w;
   wire [7:0] _00003a337_00003a_00003areg__0;
   wire [7:0] _00003a337_00003a_00003areg__1;
   wire [0:0] _00003a337_00003a_00003a_00003a275_00003a_00003aabus__r;
   wire [0:0] _00003a337_00003a_00003a_00003a276_00003a_00003aabus__w;
   wire [0:0] _00003a337_00003a_00003a_00003a277_00003a_00003aabus__r;
   wire [0:0] _00003a337_00003a_00003a_00003a278_00003a_00003aabus__w;
   reg [7:0] _00003a338_00003a_00003alv0;
   reg [7:0] _00003a338_00003a_00003alv1;
   reg [7:0] _00003a338_00003a_00003arv0;
   reg [7:0] _00003a338_00003a_00003arv1;
   reg _00003a338_00003a_00003alvok0;
   reg _00003a338_00003a_00003alvok1;
   reg _00003a338_00003a_00003arvok0;
   reg _00003a338_00003a_00003arvok1;
   reg _00003a338_00003a_00003arun;
   wire [7:0] _00003a339_00003a_00003areg__0;
   wire [7:0] _00003a339_00003a_00003areg__1;
   wire [0:0] _00003a339_00003a_00003a_00003a293_00003a_00003aabus__r;
   wire [0:0] _00003a339_00003a_00003a_00003a294_00003a_00003aabus__w;
   wire [0:0] _00003a339_00003a_00003a_00003a295_00003a_00003aabus__r;
   wire [0:0] _00003a339_00003a_00003a_00003a296_00003a_00003aabus__w;
   wire [7:0] _00005e_0000600;
   wire [7:0] _00005e_0000601;
   wire [7:0] _00005e_0000602;
   wire [7:0] _00005e_0000603;

   _____00003aT0_00003a_00003afunc0_00003aT0 func0(.z__value(_00005e_0000600),.a(_00005e_0000601));
   _____00003aT0_00003a_00003afunc1_00003aT0 func1(.z__value(_00005e_0000602),.a(_00005e_0000603));
   assign _00005e_0000600 = z0__val;

   assign a0__val = _00005e_0000601;

   assign _00005e_0000602 = z1__val;

   assign a1__val = _00005e_0000603;

   assign _00003a14 = _00003a331_00003a_00003adbus__r;

   assign _00003a12 = _00003a331_00003a_00003atrig__r;

   assign _00003a13 = _00003a331_00003a_00003aabus__r;

   assign _00003a16 = _00003a331_00003a_00003atrig__w;

   assign _00003a17 = _00003a331_00003a_00003aabus__w;

   assign _00003a18 = _00003a331_00003a_00003adbus__w;

   assign _00003a43 = _00003a332_00003a_00003adbus__r;

   assign _00003a41 = _00003a332_00003a_00003atrig__r;

   assign _00003a42 = _00003a332_00003a_00003aabus__r;

   assign _00003a45 = _00003a332_00003a_00003atrig__w;

   assign _00003a46 = _00003a332_00003a_00003aabus__w;

   assign _00003a47 = _00003a332_00003a_00003adbus__w;

   assign _00003a72 = _00003a333_00003a_00003adbus__r;

   assign _00003a70 = _00003a333_00003a_00003atrig__r;

   assign _00003a71 = _00003a333_00003a_00003aabus__r;

   assign _00003a74 = _00003a333_00003a_00003atrig__w;

   assign _00003a75 = _00003a333_00003a_00003aabus__w;

   assign _00003a76 = _00003a333_00003a_00003adbus__w;

   assign _00003a89 = _00003a334_00003a_00003areg__0;

   assign _00003a90 = _00003a334_00003a_00003areg__1;

   assign _00003a120 = _00003a336_00003a_00003areg__0;

   assign _00003a121 = _00003a336_00003a_00003areg__1;

   assign _00003a135 = _00003a336_00003a_00003areg__0;

   assign _00003a136 = _00003a336_00003a_00003areg__1;

   assign _00003a137 = _00003a336_00003a_00003a_00003a269_00003a_00003aabus__w;

   assign _00003a150 = _00003a337_00003a_00003areg__0;

   assign _00003a151 = _00003a337_00003a_00003areg__1;

   assign _00003a181 = _00003a339_00003a_00003areg__0;

   assign _00003a182 = _00003a339_00003a_00003areg__1;

   always @( posedge clk ) begin

      if (ackB) begin
         z0__val <= _00003a150;
         z1__val <= _00003a151;
         _00003a181 <= a0__val;
         _00003a182 <= a1__val;
         ack <= 32'd1;
      end

   end

   always @( posedge clk ) begin

      if ((rst == 32'd1)) begin
         _00003a137 <= 32'd0;
      end

      if ((rst == 32'd1)) begin
         _00003a75 <= -32'd1;
      end

      _00003a74 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a46 <= -32'd1;
      end

      _00003a45 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a17 <= -32'd1;
      end

      _00003a16 <= 32'd0;

      if (fill) begin
         if ((rst == 32'd0)) begin
            _00003a17 <= (_00003a17 + 32'd1);
            _00003a16 <= 32'd1;
            _00003a18 <= val;
         end
         if ((rst == 32'd0)) begin
            _00003a46 <= (_00003a46 + 32'd1);
            _00003a45 <= 32'd1;
            _00003a47 <= val;
         end
         if ((rst == 32'd0)) begin
            _00003a75 <= (_00003a75 + 32'd1);
            _00003a74 <= 32'd1;
            _00003a76 <= val;
         end
         if ((rst == 32'd0)) begin
            case(_00003a137)
               32'd0: _00003a135 <= val;
               32'd1: _00003a136 <= val;
            endcase
            _00003a137 <= (_00003a137 + 32'd1);
         end
      end

   end

   initial begin

      clk = 32'd0;

      rst = 32'd0;

      req = 32'd0;

      val = 32'd0;

      fill = 32'd0;

      #10000

      rst = 32'd1;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      rst = 32'd0;

      fill = 32'd1;

      val = 32'd1;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      #10000

      fill = 32'd0;

      clk = 32'd1;

      clk = 32'd0;

      req = 32'd1;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      if ((ackB == 32'd1)) begin
         req = 32'd0;
      end

      #10000

   end

   always @( negedge clk ) begin

      _00003a331_00003a_00003adbus__r <= _00003a331_00003a_00003amem[_00003a331_00003a_00003aabus__r];

      if (_00003a331_00003a_00003atrig__w) begin
         _00003a331_00003a_00003amem[_00003a331_00003a_00003aabus__w] <= _00003a331_00003a_00003adbus__w;
      end

   end

   always @( negedge clk ) begin

      _00003a332_00003a_00003adbus__r <= _00003a332_00003a_00003amem[_00003a332_00003a_00003aabus__r];

      if (_00003a332_00003a_00003atrig__w) begin
         _00003a332_00003a_00003amem[_00003a332_00003a_00003aabus__w] <= _00003a332_00003a_00003adbus__w;
      end

   end

   always @( negedge clk ) begin

      _00003a333_00003a_00003adbus__r <= _00003a333_00003a_00003amem[_00003a333_00003a_00003aabus__r];

      if (_00003a333_00003a_00003atrig__w) begin
         _00003a333_00003a_00003amem[_00003a333_00003a_00003aabus__w] <= _00003a333_00003a_00003adbus__w;
      end

   end

   always @( posedge clk ) begin

      if ((rst == 32'd1)) begin
         _00003a42 <= -32'd1;
      end

      _00003a41 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a13 <= -32'd1;
      end

      _00003a12 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a71 <= -32'd1;
      end

      _00003a70 <= 32'd0;

      ackA <= 32'd0;

      _00003a335_00003a_00003arun <= 32'd0;

      if ((req | _00003a335_00003a_00003arun)) begin
         _00003a335_00003a_00003arun <= 32'd1;
         if ((rst == 32'd0)) begin
            if ((_00003a70 == 32'd1)) begin
               _00003a335_00003a_00003arv <= _00003a72;
               _00003a335_00003a_00003arvok <= 32'd1;
            end
            _00003a71 <= (_00003a71 + 32'd1);
            _00003a70 <= 32'd1;
         end
         if ((rst == 32'd0)) begin
            if ((_00003a12 == 32'd1)) begin
               _00003a335_00003a_00003alv0 <= _00003a14;
               _00003a335_00003a_00003alvok0 <= 32'd1;
            end
            _00003a13 <= (_00003a13 + 32'd1);
            _00003a12 <= 32'd1;
         end
         if ((_00003a335_00003a_00003alvok0 & _00003a335_00003a_00003arvok)) begin
            ackA <= 32'd1;
            _00003a335_00003a_00003arun <= 32'd0;
            _00003a335_00003a_00003aav0 <= (_00003a335_00003a_00003aav0 + (_00003a335_00003a_00003alv0 * _00003a335_00003a_00003arv));
            _00003a89 <= ((_00003a335_00003a_00003aav0 + (_00003a335_00003a_00003alv0 * _00003a335_00003a_00003arv)) + (_00003a335_00003a_00003alv0 * _00003a335_00003a_00003arv));
         end
         if ((rst == 32'd0)) begin
            if ((_00003a41 == 32'd1)) begin
               _00003a335_00003a_00003alv1 <= _00003a43;
               _00003a335_00003a_00003alvok1 <= 32'd1;
            end
            _00003a42 <= (_00003a42 + 32'd1);
            _00003a41 <= 32'd1;
         end
         if ((_00003a335_00003a_00003alvok1 & _00003a335_00003a_00003arvok)) begin
            ackA <= 32'd1;
            _00003a335_00003a_00003arun <= 32'd0;
            _00003a335_00003a_00003aav1 <= (_00003a335_00003a_00003aav1 + (_00003a335_00003a_00003alv1 * _00003a335_00003a_00003arv));
            _00003a90 <= ((_00003a335_00003a_00003aav1 + (_00003a335_00003a_00003alv1 * _00003a335_00003a_00003arv)) + (_00003a335_00003a_00003alv1 * _00003a335_00003a_00003arv));
         end
      end
      else begin
         _00003a335_00003a_00003arvok <= 32'd0;
         _00003a335_00003a_00003alvok0 <= 32'd0;
         _00003a335_00003a_00003aav0 <= 32'd0;
         _00003a335_00003a_00003alvok1 <= 32'd0;
         _00003a335_00003a_00003aav1 <= 32'd0;
      end

   end

   always @( posedge clk ) begin

      ackB <= 32'd0;

      _00003a338_00003a_00003arun <= 32'd0;

      if ((ackA | _00003a338_00003a_00003arun)) begin
         _00003a338_00003a_00003arun <= 32'd1;
         _00003a338_00003a_00003alv0 <= _00003a89;
         _00003a338_00003a_00003alvok0 <= 32'd1;
         _00003a338_00003a_00003arv0 <= _00003a120;
         _00003a338_00003a_00003arvok0 <= 32'd1;
         if ((_00003a338_00003a_00003alvok0 & _00003a338_00003a_00003arvok0)) begin
            _00003a338_00003a_00003arun <= 32'd0;
            ackB <= 32'd1;
            _00003a150 <= (_00003a338_00003a_00003alv0 + _00003a338_00003a_00003arv0);
         end
         _00003a338_00003a_00003alv1 <= _00003a90;
         _00003a338_00003a_00003alvok1 <= 32'd1;
         _00003a338_00003a_00003arv1 <= _00003a121;
         _00003a338_00003a_00003arvok1 <= 32'd1;
         if ((_00003a338_00003a_00003alvok1 & _00003a338_00003a_00003arvok1)) begin
            _00003a338_00003a_00003arun <= 32'd0;
            ackB <= 32'd1;
            _00003a151 <= (_00003a338_00003a_00003alv1 + _00003a338_00003a_00003arv1);
         end
      end
      else begin
         _00003a338_00003a_00003alvok0 <= 32'd0;
         _00003a338_00003a_00003arvok0 <= 32'd0;
         _00003a338_00003a_00003alvok1 <= 32'd0;
         _00003a338_00003a_00003arvok1 <= 32'd0;
      end

   end

endmodule