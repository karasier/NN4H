`timescale 1ps/1ps

module _____00003aT0_00003a_00003asubtractor_00003aT0( a, b, s ); 
   input [3:0] a;
   input [3:0] b;
   output [4:0] s;

   assign s = (a - b);

endmodule