`timescale 1ps/1ps

module _____00003aT0( ); 
   reg clk;
   reg rst;
   wire [7:0] _00003a76_00003a_00003areg__0;
   wire [7:0] _00003a76_00003a_00003areg__1;
   wire [0:0] _00003a76_00003a_00003a_00003a65_00003a_00003aabus__r;
   wire [0:0] _00003a76_00003a_00003a_00003a66_00003a_00003aabus__w;
   wire [0:0] _00003a76_00003a_00003a_00003a67_00003a_00003aabus__r;
   wire [0:0] _00003a76_00003a_00003a_00003a68_00003a_00003aabus__w;
   wire [7:0] _00003a77_00003a_00003areg__0;
   wire [7:0] _00003a77_00003a_00003areg__1;
   wire [0:0] _00003a77_00003a_00003a_00003a72_00003a_00003aabus__r;
   wire [0:0] _00003a77_00003a_00003a_00003a73_00003a_00003aabus__w;
   wire [0:0] _00003a77_00003a_00003a_00003a74_00003a_00003aabus__r;
   wire [0:0] _00003a77_00003a_00003a_00003a75_00003a_00003aabus__w;
   wire _00005e_0000600;
   wire _00005e_0000601;

   _____00003aT0_00003a_00003alayer_00003aT0 layer(.clk(_00005e_0000600),.rst(_00005e_0000601));
   assign _00005e_0000600 = clk;

   assign _00005e_0000601 = rst;

   initial begin

      clk = 32'd0;

      rst = 32'd0;

   end

endmodule