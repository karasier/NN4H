`timescale 1ps/1ps

module _____00003aT0( addr, data ); 
   input [7:0] addr;
   output [255:0] data;
   reg signed[7:0] content  [255:0];

   assign data = content[addr];

   initial begin

      content[32'd0] = 53'b-1.0;

      content[32'd1] = 53'b-1.0;

      content[32'd2] = 53'b-1.0;

      content[32'd3] = 53'b-1.0;

      content[32'd4] = 53'b-1.0;

      content[32'd5] = 53'b-1.0;

      content[32'd6] = 53'b-1.0;

      content[32'd7] = 53'b-1.0;

      content[32'd8] = 53'b-1.0;

      content[32'd9] = 53'b-1.0;

      content[32'd10] = 53'b-1.0;

      content[32'd11] = 53'b-1.0;

      content[32'd12] = 53'b-1.0;

      content[32'd13] = 53'b-1.0;

      content[32'd14] = 53'b-1.0;

      content[32'd15] = 53'b-1.0;

      content[32'd16] = 53'b-1.0;

      content[32'd17] = 53'b-1.0;

      content[32'd18] = 53'b-1.0;

      content[32'd19] = 53'b-1.0;

      content[32'd20] = 53'b-1.0;

      content[32'd21] = 53'b-1.0;

      content[32'd22] = 53'b-1.0;

      content[32'd23] = 53'b-1.0;

      content[32'd24] = 53'b-1.0;

      content[32'd25] = 53'b-1.0;

      content[32'd26] = 53'b-1.0;

      content[32'd27] = 53'b-1.0;

      content[32'd28] = 53'b-1.0;

      content[32'd29] = 53'b-1.0;

      content[32'd30] = 53'b-1.0;

      content[32'd31] = 53'b-1.0;

      content[32'd32] = 53'b-1.0;

      content[32'd33] = 53'b-1.0;

      content[32'd34] = 53'b-1.0;

      content[32'd35] = 53'b-1.0;

      content[32'd36] = 53'b-1.0;

      content[32'd37] = 53'b-1.0;

      content[32'd38] = 53'b-1.0;

      content[32'd39] = 53'b-1.0;

      content[32'd40] = 53'b-1.0;

      content[32'd41] = 53'b-1.0;

      content[32'd42] = 53'b-1.0;

      content[32'd43] = 53'b-1.0;

      content[32'd44] = 53'b-1.0;

      content[32'd45] = 53'b-1.0;

      content[32'd46] = 53'b-1.0;

      content[32'd47] = 53'b-1.0;

      content[32'd48] = 53'b-1.0;

      content[32'd49] = 53'b-1.0;

      content[32'd50] = 53'b-1.0;

      content[32'd51] = 53'b-1.0;

      content[32'd52] = 53'b-1.0;

      content[32'd53] = 53'b-1.0;

      content[32'd54] = 53'b-1.0;

      content[32'd55] = 53'b-1.0;

      content[32'd56] = 53'b-1.0;

      content[32'd57] = 53'b-1.0;

      content[32'd58] = 53'b-1.0;

      content[32'd59] = 53'b-1.0;

      content[32'd60] = 53'b-1.0;

      content[32'd61] = 53'b-1.0;

      content[32'd62] = 53'b-1.0;

      content[32'd63] = 53'b-1.0;

      content[32'd64] = 53'b-1.0;

      content[32'd65] = 53'b-1.0;

      content[32'd66] = 53'b-1.0;

      content[32'd67] = 53'b-1.0;

      content[32'd68] = 53'b-1.0;

      content[32'd69] = 53'b-1.0;

      content[32'd70] = 53'b-1.0;

      content[32'd71] = 53'b-1.0;

      content[32'd72] = 53'b-1.0;

      content[32'd73] = 53'b-1.0;

      content[32'd74] = 53'b-1.0;

      content[32'd75] = 53'b-1.0;

      content[32'd76] = 53'b-1.0;

      content[32'd77] = 53'b-1.0;

      content[32'd78] = 53'b-1.0;

      content[32'd79] = 53'b-1.0;

      content[32'd80] = 53'b-1.0;

      content[32'd81] = 53'b-1.0;

      content[32'd82] = 53'b-1.0;

      content[32'd83] = 53'b-1.0;

      content[32'd84] = 53'b-1.0;

      content[32'd85] = 53'b-1.0;

      content[32'd86] = 53'b-1.0;

      content[32'd87] = 53'b-1.0;

      content[32'd88] = 53'b-1.0;

      content[32'd89] = 53'b-1.0;

      content[32'd90] = 53'b-1.0;

      content[32'd91] = 53'b-1.0;

      content[32'd92] = 53'b-1.0;

      content[32'd93] = 53'b-1.0;

      content[32'd94] = 53'b-1.0;

      content[32'd95] = 53'b-1.0;

      content[32'd96] = 53'b-1.0;

      content[32'd97] = 53'b-1.0;

      content[32'd98] = 53'b-1.0;

      content[32'd99] = 53'b-1.0;

      content[32'd100] = 53'b-1.0;

      content[32'd101] = 53'b-1.0;

      content[32'd102] = 53'b-1.0;

      content[32'd103] = 53'b-1.0;

      content[32'd104] = 53'b-1.0;

      content[32'd105] = 53'b-1.0;

      content[32'd106] = 53'b-1.0;

      content[32'd107] = 53'b-1.0;

      content[32'd108] = 53'b-1.0;

      content[32'd109] = 53'b-0.9999999999999999;

      content[32'd110] = 53'b-0.9999999999999996;

      content[32'd111] = 53'b-0.9999999999999966;

      content[32'd112] = 53'b-0.9999999999999747;

      content[32'd113] = 53'b-0.9999999999998128;

      content[32'd114] = 53'b-0.9999999999986171;

      content[32'd115] = 53'b-0.9999999999897818;

      content[32'd116] = 53'b-0.9999999999244973;

      content[32'd117] = 53'b-0.9999999994421064;

      content[32'd118] = 53'b-0.9999999958776927;

      content[32'd119] = 53'b-0.999999969540041;

      content[32'd120] = 53'b-0.9999997749296758;

      content[32'd121] = 53'b-0.9999983369439447;

      content[32'd122] = 53'b-0.9999877116507956;

      content[32'd123] = 53'b-0.9999092042625951;

      content[32'd124] = 53'b-0.999329299739067;

      content[32'd125] = 53'b-0.9950547536867305;

      content[32'd126] = 53'b-0.9640275800758169;

      content[32'd127] = 53'b-0.7615941559557649;

      content[32'd128] = 53'b0.0;

      content[32'd129] = 53'b0.7615941559557649;

      content[32'd130] = 53'b0.9640275800758169;

      content[32'd131] = 53'b0.9950547536867305;

      content[32'd132] = 53'b0.999329299739067;

      content[32'd133] = 53'b0.9999092042625951;

      content[32'd134] = 53'b0.9999877116507956;

      content[32'd135] = 53'b0.9999983369439447;

      content[32'd136] = 53'b0.9999997749296758;

      content[32'd137] = 53'b0.999999969540041;

      content[32'd138] = 53'b0.9999999958776927;

      content[32'd139] = 53'b0.9999999994421064;

      content[32'd140] = 53'b0.9999999999244973;

      content[32'd141] = 53'b0.9999999999897818;

      content[32'd142] = 53'b0.9999999999986171;

      content[32'd143] = 53'b0.9999999999998128;

      content[32'd144] = 53'b0.9999999999999747;

      content[32'd145] = 53'b0.9999999999999966;

      content[32'd146] = 53'b0.9999999999999996;

      content[32'd147] = 53'b0.9999999999999999;

      content[32'd148] = 53'b1.0;

      content[32'd149] = 53'b1.0;

      content[32'd150] = 53'b1.0;

      content[32'd151] = 53'b1.0;

      content[32'd152] = 53'b1.0;

      content[32'd153] = 53'b1.0;

      content[32'd154] = 53'b1.0;

      content[32'd155] = 53'b1.0;

      content[32'd156] = 53'b1.0;

      content[32'd157] = 53'b1.0;

      content[32'd158] = 53'b1.0;

      content[32'd159] = 53'b1.0;

      content[32'd160] = 53'b1.0;

      content[32'd161] = 53'b1.0;

      content[32'd162] = 53'b1.0;

      content[32'd163] = 53'b1.0;

      content[32'd164] = 53'b1.0;

      content[32'd165] = 53'b1.0;

      content[32'd166] = 53'b1.0;

      content[32'd167] = 53'b1.0;

      content[32'd168] = 53'b1.0;

      content[32'd169] = 53'b1.0;

      content[32'd170] = 53'b1.0;

      content[32'd171] = 53'b1.0;

      content[32'd172] = 53'b1.0;

      content[32'd173] = 53'b1.0;

      content[32'd174] = 53'b1.0;

      content[32'd175] = 53'b1.0;

      content[32'd176] = 53'b1.0;

      content[32'd177] = 53'b1.0;

      content[32'd178] = 53'b1.0;

      content[32'd179] = 53'b1.0;

      content[32'd180] = 53'b1.0;

      content[32'd181] = 53'b1.0;

      content[32'd182] = 53'b1.0;

      content[32'd183] = 53'b1.0;

      content[32'd184] = 53'b1.0;

      content[32'd185] = 53'b1.0;

      content[32'd186] = 53'b1.0;

      content[32'd187] = 53'b1.0;

      content[32'd188] = 53'b1.0;

      content[32'd189] = 53'b1.0;

      content[32'd190] = 53'b1.0;

      content[32'd191] = 53'b1.0;

      content[32'd192] = 53'b1.0;

      content[32'd193] = 53'b1.0;

      content[32'd194] = 53'b1.0;

      content[32'd195] = 53'b1.0;

      content[32'd196] = 53'b1.0;

      content[32'd197] = 53'b1.0;

      content[32'd198] = 53'b1.0;

      content[32'd199] = 53'b1.0;

      content[32'd200] = 53'b1.0;

      content[32'd201] = 53'b1.0;

      content[32'd202] = 53'b1.0;

      content[32'd203] = 53'b1.0;

      content[32'd204] = 53'b1.0;

      content[32'd205] = 53'b1.0;

      content[32'd206] = 53'b1.0;

      content[32'd207] = 53'b1.0;

      content[32'd208] = 53'b1.0;

      content[32'd209] = 53'b1.0;

      content[32'd210] = 53'b1.0;

      content[32'd211] = 53'b1.0;

      content[32'd212] = 53'b1.0;

      content[32'd213] = 53'b1.0;

      content[32'd214] = 53'b1.0;

      content[32'd215] = 53'b1.0;

      content[32'd216] = 53'b1.0;

      content[32'd217] = 53'b1.0;

      content[32'd218] = 53'b1.0;

      content[32'd219] = 53'b1.0;

      content[32'd220] = 53'b1.0;

      content[32'd221] = 53'b1.0;

      content[32'd222] = 53'b1.0;

      content[32'd223] = 53'b1.0;

      content[32'd224] = 53'b1.0;

      content[32'd225] = 53'b1.0;

      content[32'd226] = 53'b1.0;

      content[32'd227] = 53'b1.0;

      content[32'd228] = 53'b1.0;

      content[32'd229] = 53'b1.0;

      content[32'd230] = 53'b1.0;

      content[32'd231] = 53'b1.0;

      content[32'd232] = 53'b1.0;

      content[32'd233] = 53'b1.0;

      content[32'd234] = 53'b1.0;

      content[32'd235] = 53'b1.0;

      content[32'd236] = 53'b1.0;

      content[32'd237] = 53'b1.0;

      content[32'd238] = 53'b1.0;

      content[32'd239] = 53'b1.0;

      content[32'd240] = 53'b1.0;

      content[32'd241] = 53'b1.0;

      content[32'd242] = 53'b1.0;

      content[32'd243] = 53'b1.0;

      content[32'd244] = 53'b1.0;

      content[32'd245] = 53'b1.0;

      content[32'd246] = 53'b1.0;

      content[32'd247] = 53'b1.0;

      content[32'd248] = 53'b1.0;

      content[32'd249] = 53'b1.0;

      content[32'd250] = 53'b1.0;

      content[32'd251] = 53'b1.0;

      content[32'd252] = 53'b1.0;

      content[32'd253] = 53'b1.0;

      content[32'd254] = 53'b1.0;

      content[32'd255] = 53'b1.0;

      content[32'd256] = 53'b1.0;

   end

endmodule