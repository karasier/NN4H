`timescale 1ps/1ps

module _____00003aT0_00003a_00003alayer_00003aT0( clk,   input clk;
   input rst;
   wire req;

endmodule