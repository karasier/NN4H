`timescale 1ps/1ps

module _____00003aT0( ); 

   _____00003aT0_00003a_00003aadder_00003aT0 adder);
   _____00003aT0_00003a_00003asubtractor_00003aT0 subtractor);
   _____00003aT0_00003a_00003amultiplier_00003aT0 multiplier);
   _____00003aT0_00003a_00003adivider_00003aT0 divider);
endmodule