`timescale 1ps/1ps

module _____00003aT0_00003a_00003atanh__neural__network_00003aT0_00003a_00003alayer1_00003aT00_00003a_00003afunc0_00003aT20( z__value, a ); 
   input signed[7:0] z__value;
   output signed[7:0] a;
   wire signed[7:0] base;
   wire signed[7:0] next__data;
   wire [3:0] address;
   wire signed[7:0] remaining;
   wire signed[7:0] change;
   wire [3:0] _00005e_000060605;
   wire signed[7:0] _00005e_000060606;
   wire signed[7:0] _00005e_000060607;
   wire signed[7:0] _00005e_000060608;
   wire signed[7:0] _00005e_000060609;
   wire signed[7:0] _00005e_000060610;
   wire signed[7:0] _00005e_000060611;
   wire signed[7:0] _00005e_000060612;

   _____00003aT0_00003a_00003atanh__neural__network_00003aT0_00003a_00003alayer1_00003aT00_00003a_00003afunc0_00003aT20_00003a_00003amy__lut_00003aT40 my__lut(.address(_00005e_000060605),.base(_00005e_000060606),.next__data(_00005e_000060607));
   _____00003aT0_00003a_00003atanh__neural__network_00003aT0_00003a_00003alayer1_00003aT00_00003a_00003afunc0_00003aT20_00003a_00003amy__interpolator_00003aT40 my__interpolator(.base(_00005e_000060608),.next__data(_00005e_000060609),.change(_00005e_000060610),.remaining(_00005e_000060611),.interpolated__value(_00005e_000060612));
   assign address = z__value[7:4];

   assign remaining = {{1'b0,1'b0,1'b0,1'b0},z__value[3:0]};

   assign change = {{1'b0,1'b0,1'b0},1'b1,{1'b0,1'b0,1'b0,1'b0}};

   assign _00005e_000060605 = address;

   assign base = _00005e_000060606;

   assign next__data = _00005e_000060607;

   assign _00005e_000060608 = base;

   assign _00005e_000060609 = next__data;

   assign _00005e_000060610 = change;

   assign _00005e_000060611 = remaining;

   assign a = _00005e_000060612;

endmodule