`timescale 1ps/1ps

module _____00003aT0( ); 
   reg clk;
   reg rst;
   reg req;
   wire [7:0] _00003a14;
   reg _00003a12;
   reg [0:0] _00003a13;
   wire [7:0] _00003a43;
   reg _00003a41;
   reg [0:0] _00003a42;
   wire [7:0] _00003a72;
   reg _00003a70;
   reg [0:0] _00003a71;
   reg [7:0] _00003a89;
   reg [7:0] _00003a90;
   reg ack0;
   reg _00003a16;
   reg [0:0] _00003a17;
   reg [7:0] _00003a18;
   reg _00003a45;
   reg [0:0] _00003a46;
   reg [7:0] _00003a47;
   reg _00003a74;
   reg [0:0] _00003a75;
   reg [7:0] _00003a76;
   reg [7:0] val;
   wire _00003a185_00003a_00003atrig__r;
   wire _00003a185_00003a_00003atrig__w;
   reg [7:0] _00003a185_00003a_00003adbus__r;
   wire [7:0] _00003a185_00003a_00003adbus__w;
   wire [0:0] _00003a185_00003a_00003aabus__r;
   wire [0:0] _00003a185_00003a_00003aabus__w;
   reg [7:0] _00003a185_00003a_00003amem  [0:1];
   wire _00003a186_00003a_00003atrig__r;
   wire _00003a186_00003a_00003atrig__w;
   reg [7:0] _00003a186_00003a_00003adbus__r;
   wire [7:0] _00003a186_00003a_00003adbus__w;
   wire [0:0] _00003a186_00003a_00003aabus__r;
   wire [0:0] _00003a186_00003a_00003aabus__w;
   reg [7:0] _00003a186_00003a_00003amem  [0:1];
   wire _00003a187_00003a_00003atrig__r;
   wire _00003a187_00003a_00003atrig__w;
   reg [7:0] _00003a187_00003a_00003adbus__r;
   wire [7:0] _00003a187_00003a_00003adbus__w;
   wire [0:0] _00003a187_00003a_00003aabus__r;
   wire [0:0] _00003a187_00003a_00003aabus__w;
   reg [7:0] _00003a187_00003a_00003amem  [0:1];
   wire [7:0] _00003a188_00003a_00003areg__0;
   wire [7:0] _00003a188_00003a_00003areg__1;
   wire [0:0] _00003a188_00003a_00003a_00003a145_00003a_00003aabus__r;
   wire [0:0] _00003a188_00003a_00003a_00003a146_00003a_00003aabus__w;
   wire [0:0] _00003a188_00003a_00003a_00003a147_00003a_00003aabus__r;
   wire [0:0] _00003a188_00003a_00003a_00003a148_00003a_00003aabus__w;
   reg [7:0] _00003a189_00003a_00003alv0;
   reg [7:0] _00003a189_00003a_00003alv1;
   reg [7:0] _00003a189_00003a_00003aav0;
   reg [7:0] _00003a189_00003a_00003aav1;
   reg [7:0] _00003a189_00003a_00003arv;
   reg _00003a189_00003a_00003alvok0;
   reg _00003a189_00003a_00003alvok1;
   reg _00003a189_00003a_00003arvok;
   reg _00003a189_00003a_00003arun;

   assign _00003a14 = _00003a185_00003a_00003adbus__r;

   assign _00003a12 = _00003a185_00003a_00003atrig__r;

   assign _00003a13 = _00003a185_00003a_00003aabus__r;

   assign _00003a16 = _00003a185_00003a_00003atrig__w;

   assign _00003a17 = _00003a185_00003a_00003aabus__w;

   assign _00003a18 = _00003a185_00003a_00003adbus__w;

   assign _00003a43 = _00003a186_00003a_00003adbus__r;

   assign _00003a41 = _00003a186_00003a_00003atrig__r;

   assign _00003a42 = _00003a186_00003a_00003aabus__r;

   assign _00003a45 = _00003a186_00003a_00003atrig__w;

   assign _00003a46 = _00003a186_00003a_00003aabus__w;

   assign _00003a47 = _00003a186_00003a_00003adbus__w;

   assign _00003a72 = _00003a187_00003a_00003adbus__r;

   assign _00003a70 = _00003a187_00003a_00003atrig__r;

   assign _00003a71 = _00003a187_00003a_00003aabus__r;

   assign _00003a74 = _00003a187_00003a_00003atrig__w;

   assign _00003a75 = _00003a187_00003a_00003aabus__w;

   assign _00003a76 = _00003a187_00003a_00003adbus__w;

   assign _00003a89 = _00003a188_00003a_00003areg__0;

   assign _00003a90 = _00003a188_00003a_00003areg__1;

   always @( posedge clk ) begin

      if ((rst == 32'd1)) begin
         _00003a75 <= -32'd1;
      end

      _00003a74 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a46 <= -32'd1;
      end

      _00003a45 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a17 <= -32'd1;
      end

      _00003a16 <= 32'd0;

      if ((rst == 32'd0)) begin
         _00003a17 <= (_00003a17 + 32'd1);
         _00003a16 <= 32'd1;
         _00003a18 <= val;
      end

      if ((rst == 32'd0)) begin
         _00003a46 <= (_00003a46 + 32'd1);
         _00003a45 <= 32'd1;
         _00003a47 <= (val + 32'd1);
      end

      if ((rst == 32'd0)) begin
         _00003a75 <= (_00003a75 + 32'd1);
         _00003a74 <= 32'd1;
         _00003a76 <= (val + 32'd1);
      end

   end

   initial begin

      req = 32'd0;

      clk = 32'd0;

      rst = 32'd0;

      val = 32'd0;

      #10000

      rst = 32'd1;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      rst = 32'd0;

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      val = (val + 32'd1);

      #10000

      clk = 32'd1;

      #10000

      clk = 32'd0;

      val = (val + 32'd1);

      #10000

   end

   always @( negedge clk ) begin

      _00003a185_00003a_00003adbus__r <= _00003a185_00003a_00003amem[_00003a185_00003a_00003aabus__r];

      if (_00003a185_00003a_00003atrig__w) begin
         _00003a185_00003a_00003amem[_00003a185_00003a_00003aabus__w] <= _00003a185_00003a_00003adbus__w;
      end

   end

   always @( negedge clk ) begin

      _00003a186_00003a_00003adbus__r <= _00003a186_00003a_00003amem[_00003a186_00003a_00003aabus__r];

      if (_00003a186_00003a_00003atrig__w) begin
         _00003a186_00003a_00003amem[_00003a186_00003a_00003aabus__w] <= _00003a186_00003a_00003adbus__w;
      end

   end

   always @( negedge clk ) begin

      _00003a187_00003a_00003adbus__r <= _00003a187_00003a_00003amem[_00003a187_00003a_00003aabus__r];

      if (_00003a187_00003a_00003atrig__w) begin
         _00003a187_00003a_00003amem[_00003a187_00003a_00003aabus__w] <= _00003a187_00003a_00003adbus__w;
      end

   end

   always @( posedge clk ) begin

      if ((rst == 32'd1)) begin
         _00003a42 <= -32'd1;
      end

      _00003a41 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a13 <= -32'd1;
      end

      _00003a12 <= 32'd0;

      if ((rst == 32'd1)) begin
         _00003a71 <= -32'd1;
      end

      _00003a70 <= 32'd0;

      ack0 <= 32'd0;

      _00003a189_00003a_00003arun <= 32'd0;

      if ((req | _00003a189_00003a_00003arun)) begin
         _00003a189_00003a_00003arun <= 32'd1;
         if ((rst == 32'd0)) begin
            if ((_00003a70 == 32'd1)) begin
               _00003a189_00003a_00003arv <= _00003a72;
               _00003a189_00003a_00003arvok <= 32'd1;
            end
            _00003a71 <= (_00003a71 + 32'd1);
            _00003a70 <= 32'd1;
         end
         if ((rst == 32'd0)) begin
            if ((_00003a12 == 32'd1)) begin
               _00003a189_00003a_00003alv0 <= _00003a14;
               _00003a189_00003a_00003alvok0 <= 32'd1;
            end
            _00003a13 <= (_00003a13 + 32'd1);
            _00003a12 <= 32'd1;
         end
         if ((_00003a189_00003a_00003alvok0 & _00003a189_00003a_00003arvok)) begin
            ack0 <= 32'd1;
            _00003a189_00003a_00003arun <= 32'd0;
            _00003a189_00003a_00003aav0 <= (_00003a189_00003a_00003aav0 + (_00003a189_00003a_00003alv0 * _00003a189_00003a_00003arv));
            _00003a89 <= ((_00003a189_00003a_00003aav0 + (_00003a189_00003a_00003alv0 * _00003a189_00003a_00003arv)) + (_00003a189_00003a_00003alv0 * _00003a189_00003a_00003arv));
         end
         if ((rst == 32'd0)) begin
            if ((_00003a41 == 32'd1)) begin
               _00003a189_00003a_00003alv1 <= _00003a43;
               _00003a189_00003a_00003alvok1 <= 32'd1;
            end
            _00003a42 <= (_00003a42 + 32'd1);
            _00003a41 <= 32'd1;
         end
         if ((_00003a189_00003a_00003alvok1 & _00003a189_00003a_00003arvok)) begin
            ack0 <= 32'd1;
            _00003a189_00003a_00003arun <= 32'd0;
            _00003a189_00003a_00003aav1 <= (_00003a189_00003a_00003aav1 + (_00003a189_00003a_00003alv1 * _00003a189_00003a_00003arv));
            _00003a90 <= ((_00003a189_00003a_00003aav1 + (_00003a189_00003a_00003alv1 * _00003a189_00003a_00003arv)) + (_00003a189_00003a_00003alv1 * _00003a189_00003a_00003arv));
         end
      end
      else begin
         _00003a189_00003a_00003arvok <= 32'd0;
         _00003a189_00003a_00003alvok0 <= 32'd0;
         _00003a189_00003a_00003aav0 <= 32'd0;
         _00003a189_00003a_00003alvok1 <= 32'd0;
         _00003a189_00003a_00003aav1 <= 32'd0;
      end

   end

endmodule