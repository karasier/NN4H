`timescale 1ps/1ps

module _____00003aT0_00003a_00003atanh_00003aT0_00003a_00003amy__table_00003aT0( addr, base, next__data ); 
   input [7:0] addr;
   output [31:0] base;
   output reg [31:0] next__data;
   reg [31:0] lut  [0:255];

   assign base = lut[addr];

   always @( * ) begin

      if ((addr == 32'd255)) begin
         next__data <= lut[addr];
      end
      else begin
         next__data <= lut[(addr + 32'd1)];
      end

   end

   initial begin

      lut[32'd0] = 32'b00000000000000000000000000000000;

      lut[32'd1] = 32'b00000000001011111111111101110000;

      lut[32'd2] = 32'b00000000010111111111101110000000;

      lut[32'd3] = 32'b00000000100011111111000011010001;

      lut[32'd4] = 32'b00000000101111111101110000001000;

      lut[32'd5] = 32'b00000000111011111011100111001000;

      lut[32'd6] = 32'b00000001000111111000011010111101;

      lut[32'd7] = 32'b00000001010011110011111110010100;

      lut[32'd8] = 32'b00000001011111101110000100000010;

      lut[32'd9] = 32'b00000001101011100110011111000000;

      lut[32'd10] = 32'b00000001110111011101000010010010;

      lut[32'd11] = 32'b00000010000011010001100001000001;

      lut[32'd12] = 32'b00000010001111000011101110100000;

      lut[32'd13] = 32'b00000010011010110011011110001101;

      lut[32'd14] = 32'b00000010100110100000100011110000;

      lut[32'd15] = 32'b00000010110010001010110010111100;

      lut[32'd16] = 32'b00000010111101110001111111110010;

      lut[32'd17] = 32'b00000011001001010101111110011101;

      lut[32'd18] = 32'b00000011010100110110100011011010;

      lut[32'd19] = 32'b00000011100000010011100011010001;

      lut[32'd20] = 32'b00000011101011101100110010111001;

      lut[32'd21] = 32'b00000011110111000010000111011100;

      lut[32'd22] = 32'b00000100000010010011010110010010;

      lut[32'd23] = 32'b00000100001101100000010101000010;

      lut[32'd24] = 32'b00000100011000101000111001100111;

      lut[32'd25] = 32'b00000100100011101100111010001110;

      lut[32'd26] = 32'b00000100101110101100001101010100;

      lut[32'd27] = 32'b00000100111001100110101001101010;

      lut[32'd28] = 32'b00000101000100011100000110010100;

      lut[32'd29] = 32'b00000101001111001100011010101000;

      lut[32'd30] = 32'b00000101011001110111011110010011;

      lut[32'd31] = 32'b00000101100100011101001001010010;

      lut[32'd32] = 32'b00000101101110111101010011110111;

      lut[32'd33] = 32'b00000101111001010111110110101010;

      lut[32'd34] = 32'b00000110000011101100101010100111;

      lut[32'd35] = 32'b00000110001101111011101000111100;

      lut[32'd36] = 32'b00000110011000000100101011001110;

      lut[32'd37] = 32'b00000110100010000111101011010111;

      lut[32'd38] = 32'b00000110101100000100100011100100;

      lut[32'd39] = 32'b00000110110101111011001110011001;

      lut[32'd40] = 32'b00000110111111101011100110101010;

      lut[32'd41] = 32'b00000111001001010101100111100110;

      lut[32'd42] = 32'b00000111010010111001001100101011;

      lut[32'd43] = 32'b00000111011100010110010001101101;

      lut[32'd44] = 32'b00000111100101101100110010110111;

      lut[32'd45] = 32'b00000111101110111100101100100010;

      lut[32'd46] = 32'b00000111111000000101111011100001;

      lut[32'd47] = 32'b00001000000001001000011100110110;

      lut[32'd48] = 32'b00001000001010000100001101111001;

      lut[32'd49] = 32'b00001000010010111001001100010011;

      lut[32'd50] = 32'b00001000011011100111010110000000;

      lut[32'd51] = 32'b00001000100100001110101001001111;

      lut[32'd52] = 32'b00001000101100101111000100100010;

      lut[32'd53] = 32'b00001000110101001000100110101010;

      lut[32'd54] = 32'b00001000111101011011001110101011;

      lut[32'd55] = 32'b00001001000101100110111011111010;

      lut[32'd56] = 32'b00001001001101101011101101111011;

      lut[32'd57] = 32'b00001001010101101001100100100100;

      lut[32'd58] = 32'b00001001011101100000011111111001;

      lut[32'd59] = 32'b00001001100101010000100000001111;

      lut[32'd60] = 32'b00001001101100111001100110001000;

      lut[32'd61] = 32'b00001001110100011011110010010101;

      lut[32'd62] = 32'b00001001111011110111000101110110;

      lut[32'd63] = 32'b00001010000011001011100001110111;

      lut[32'd64] = 32'b00001010001010011001000111110010;

      lut[32'd65] = 32'b00001010010001011111111001001101;

      lut[32'd66] = 32'b00001010011000011111110111111010;

      lut[32'd67] = 32'b00001010011111011001000101110111;

      lut[32'd68] = 32'b00001010100110001011100101001110;

      lut[32'd69] = 32'b00001010101100110111011000010010;

      lut[32'd70] = 32'b00001010110011011100100001100001;

      lut[32'd71] = 32'b00001010111001111011000011100100;

      lut[32'd72] = 32'b00001011000000010011000001001101;

      lut[32'd73] = 32'b00001011000110100100011101010101;

      lut[32'd74] = 32'b00001011001100101111011011000000;

      lut[32'd75] = 32'b00001011010010110011111101011000;

      lut[32'd76] = 32'b00001011011000110010000111110001;

      lut[32'd77] = 32'b00001011011110101001111101100101;

      lut[32'd78] = 32'b00001011100100011011100010010100;

      lut[32'd79] = 32'b00001011101010000110111001100101;

      lut[32'd80] = 32'b00001011101111101100000111000111;

      lut[32'd81] = 32'b00001011110101001011001110101011;

      lut[32'd82] = 32'b00001011111010100100010100001010;

      lut[32'd83] = 32'b00001011111111110111011011100010;

      lut[32'd84] = 32'b00001100000101000100101000110011;

      lut[32'd85] = 32'b00001100001010001100000000000011;

      lut[32'd86] = 32'b00001100001111001101100101011101;

      lut[32'd87] = 32'b00001100010100001001011101001101;

      lut[32'd88] = 32'b00001100011000111111101011100011;

      lut[32'd89] = 32'b00001100011101110000010100110010;

      lut[32'd90] = 32'b00001100100010011011011101010001;

      lut[32'd91] = 32'b00001100100111000001001001010110;

      lut[32'd92] = 32'b00001100101011100001011101011100;

      lut[32'd93] = 32'b00001100101111111100011101111101;

      lut[32'd94] = 32'b00001100110100010010001111010111;

      lut[32'd95] = 32'b00001100111000100010110110001000;

      lut[32'd96] = 32'b00001100111100101110010110101101;

      lut[32'd97] = 32'b00001101000000110100110101101000;

      lut[32'd98] = 32'b00001101000100110110010111010110;

      lut[32'd99] = 32'b00001101001000110011000000011010;

      lut[32'd100] = 32'b00001101001100101010110101010001;

      lut[32'd101] = 32'b00001101010000011101111010011101;

      lut[32'd102] = 32'b00001101010100001100010100011011;

      lut[32'd103] = 32'b00001101010111110110000111101100;

      lut[32'd104] = 32'b00001101011011011011011000101100;

      lut[32'd105] = 32'b00001101011110111100001011111001;

      lut[32'd106] = 32'b00001101100010011000100101101101;

      lut[32'd107] = 32'b00001101100101110000101010100101;

      lut[32'd108] = 32'b00001101101001000100011110111000;

      lut[32'd109] = 32'b00001101101100010100000110111110;

      lut[32'd110] = 32'b00001101101111011111100111001101;

      lut[32'd111] = 32'b00001101110010100111000011111000;

      lut[32'd112] = 32'b00001101110101101010100001010010;

      lut[32'd113] = 32'b00001101111000101010000011101010;

      lut[32'd114] = 32'b00001101111011100101101111001110;

      lut[32'd115] = 32'b00001101111110011101101000001010;

      lut[32'd116] = 32'b00001110000001010001110010100111;

      lut[32'd117] = 32'b00001110000100000010010010101011;

      lut[32'd118] = 32'b00001110000110101111001100011010;

      lut[32'd119] = 32'b00001110001001011000100011110111;

      lut[32'd120] = 32'b00001110001011111110011101000000;

      lut[32'd121] = 32'b00001110001110100000111011110010;

      lut[32'd122] = 32'b00001110010001000000000100000110;

      lut[32'd123] = 32'b00001110010011011011111001110011;

      lut[32'd124] = 32'b00001110010101110100100000101101;

      lut[32'd125] = 32'b00001110011000001001111100100100;

      lut[32'd126] = 32'b00001110011010011100010001001000;

      lut[32'd127] = 32'b00001110011100101011100010000010;

      lut[32'd128] = 32'b00001110011110110111110010111100;

      lut[32'd129] = 32'b00001110100001000001000111011010;

      lut[32'd130] = 32'b00001110100011000111100010111110;

      lut[32'd131] = 32'b00001110100101001011001001001000;

      lut[32'd132] = 32'b00001110100111001011111101010100;

      lut[32'd133] = 32'b00001110101001001010000010111001;

      lut[32'd134] = 32'b00001110101011000101011101001111;

      lut[32'd135] = 32'b00001110101100111110001111101000;

      lut[32'd136] = 32'b00001110101110110100011101010100;

      lut[32'd137] = 32'b00001110110000101000001001011111;

      lut[32'd138] = 32'b00001110110010011001010111010010;

      lut[32'd139] = 32'b00001110110100001000001001110100;

      lut[32'd140] = 32'b00001110110101110100100100001001;

      lut[32'd141] = 32'b00001110110111011110101001010001;

      lut[32'd142] = 32'b00001110111001000110011100001000;

      lut[32'd143] = 32'b00001110111010101011111111101001;

      lut[32'd144] = 32'b00001110111100001111010110101100;

      lut[32'd145] = 32'b00001110111101110000100100000100;

      lut[32'd146] = 32'b00001110111111001111101010100011;

      lut[32'd147] = 32'b00001111000000101100101100110111;

      lut[32'd148] = 32'b00001111000010000111101101101011;

      lut[32'd149] = 32'b00001111000011100000101111100111;

      lut[32'd150] = 32'b00001111000100110111110101010001;

      lut[32'd151] = 32'b00001111000110001101000001001100;

      lut[32'd152] = 32'b00001111000111100000010101111000;

      lut[32'd153] = 32'b00001111001000110001110101110001;

      lut[32'd154] = 32'b00001111001010000001100011010001;

      lut[32'd155] = 32'b00001111001011001111100000110001;

      lut[32'd156] = 32'b00001111001100011011110000100100;

      lut[32'd157] = 32'b00001111001101100110010100111101;

      lut[32'd158] = 32'b00001111001110101111010000001011;

      lut[32'd159] = 32'b00001111001111110110100100011010;

      lut[32'd160] = 32'b00001111010000111100010011110110;

      lut[32'd161] = 32'b00001111010010000000100000100101;

      lut[32'd162] = 32'b00001111010011000011001100101101;

      lut[32'd163] = 32'b00001111010100000100011010001111;

      lut[32'd164] = 32'b00001111010101000100001011001100;

      lut[32'd165] = 32'b00001111010110000010100001100010;

      lut[32'd166] = 32'b00001111010110111111011111001100;

      lut[32'd167] = 32'b00001111010111111011000110000011;

      lut[32'd168] = 32'b00001111011000110101010111111100;

      lut[32'd169] = 32'b00001111011001101110010110101101;

      lut[32'd170] = 32'b00001111011010100110000100001000;

      lut[32'd171] = 32'b00001111011011011100100001111011;

      lut[32'd172] = 32'b00001111011100010001110001110101;

      lut[32'd173] = 32'b00001111011101000101110101100000;

      lut[32'd174] = 32'b00001111011101111000101110100111;

      lut[32'd175] = 32'b00001111011110101010011110110000;

      lut[32'd176] = 32'b00001111011111011011000111100000;

      lut[32'd177] = 32'b00001111100000001010101010011011;

      lut[32'd178] = 32'b00001111100000111001001001000001;

      lut[32'd179] = 32'b00001111100001100110100100110001;

      lut[32'd180] = 32'b00001111100010010010111111001001;

      lut[32'd181] = 32'b00001111100010111110011001100100;

      lut[32'd182] = 32'b00001111100011101000110101011100;

      lut[32'd183] = 32'b00001111100100010010010100000111;

      lut[32'd184] = 32'b00001111100100111010110110111011;

      lut[32'd185] = 32'b00001111100101100010011111001101;

      lut[32'd186] = 32'b00001111100110001001001110001111;

      lut[32'd187] = 32'b00001111100110101111000101010010;

      lut[32'd188] = 32'b00001111100111010100000101100100;

      lut[32'd189] = 32'b00001111100111111000010000010010;

      lut[32'd190] = 32'b00001111101000011011100110101001;

      lut[32'd191] = 32'b00001111101000111110001001110010;

      lut[32'd192] = 32'b00001111101001011111111010110110;

      lut[32'd193] = 32'b00001111101010000000111010111011;

      lut[32'd194] = 32'b00001111101010100001001011001000;

      lut[32'd195] = 32'b00001111101011000000101100011111;

      lut[32'd196] = 32'b00001111101011011111100000000101;

      lut[32'd197] = 32'b00001111101011111101100110111001;

      lut[32'd198] = 32'b00001111101100011011000001111100;

      lut[32'd199] = 32'b00001111101100110111110010001100;

      lut[32'd200] = 32'b00001111101101010011111000100110;

      lut[32'd201] = 32'b00001111101101101111010110000110;

      lut[32'd202] = 32'b00001111101110001010001011100111;

      lut[32'd203] = 32'b00001111101110100100011010000000;

      lut[32'd204] = 32'b00001111101110111110000010001100;

      lut[32'd205] = 32'b00001111101111010111000101000000;

      lut[32'd206] = 32'b00001111101111101111100011010001;

      lut[32'd207] = 32'b00001111110000000111011101110101;

      lut[32'd208] = 32'b00001111110000011110110101011111;

      lut[32'd209] = 32'b00001111110000110101101011000001;

      lut[32'd210] = 32'b00001111110001001011111111001011;

      lut[32'd211] = 32'b00001111110001100001110010101110;

      lut[32'd212] = 32'b00001111110001110111000110011010;

      lut[32'd213] = 32'b00001111110010001011111010111011;

      lut[32'd214] = 32'b00001111110010100000010000111111;

      lut[32'd215] = 32'b00001111110010110100001001010010;

      lut[32'd216] = 32'b00001111110011000111100100011110;

      lut[32'd217] = 32'b00001111110011011010100011001110;

      lut[32'd218] = 32'b00001111110011101101000110001100;

      lut[32'd219] = 32'b00001111110011111111001101111110;

      lut[32'd220] = 32'b00001111110100010000111011001101;

      lut[32'd221] = 32'b00001111110100100010001110011111;

      lut[32'd222] = 32'b00001111110100110011001000011001;

      lut[32'd223] = 32'b00001111110101000011101001100001;

      lut[32'd224] = 32'b00001111110101010011110010011010;

      lut[32'd225] = 32'b00001111110101100011100011100111;

      lut[32'd226] = 32'b00001111110101110010111101101100;

      lut[32'd227] = 32'b00001111110110000010000001001001;

      lut[32'd228] = 32'b00001111110110010000101110011111;

      lut[32'd229] = 32'b00001111110110011111000110001111;

      lut[32'd230] = 32'b00001111110110101101001000111000;

      lut[32'd231] = 32'b00001111110110111010110110111000;

      lut[32'd232] = 32'b00001111110111001000010000101110;

      lut[32'd233] = 32'b00001111110111010101010110110111;

      lut[32'd234] = 32'b00001111110111100010001001110000;

      lut[32'd235] = 32'b00001111110111101110101001110101;

      lut[32'd236] = 32'b00001111110111111010110111100001;

      lut[32'd237] = 32'b00001111111000000110110011010000;

      lut[32'd238] = 32'b00001111111000010010011101011010;

      lut[32'd239] = 32'b00001111111000011101110110011011;

      lut[32'd240] = 32'b00001111111000101000111110101011;

      lut[32'd241] = 32'b00001111111000110011110110100010;

      lut[32'd242] = 32'b00001111111000111110011110011001;

      lut[32'd243] = 32'b00001111111001001000110110100111;

      lut[32'd244] = 32'b00001111111001010010111111100010;

      lut[32'd245] = 32'b00001111111001011100111001100010;

      lut[32'd246] = 32'b00001111111001100110100100111011;

      lut[32'd247] = 32'b00001111111001110000000010000100;

      lut[32'd248] = 32'b00001111111001111001010001010010;

      lut[32'd249] = 32'b00001111111010000010010010111000;

      lut[32'd250] = 32'b00001111111010001011000111001010;

      lut[32'd251] = 32'b00001111111010010011101110011101;

      lut[32'd252] = 32'b00001111111010011100001001000011;

      lut[32'd253] = 32'b00001111111010100100010111001110;

      lut[32'd254] = 32'b00001111111010101100011001010010;

      lut[32'd255] = 32'b00001111111010110100001111011111;

   end

endmodule