`timescale 1ps/1ps

module _____00003aT0_00003a_00003amy__layer_00003aT0( clk, rst, req, flag, ack ); 
   input clk;
   input rst;
   input req;
   input flag;
   output reg ack;
   wire [7:0] _00003a62;
   wire [7:0] _00003a63;
   wire [7:0] _00003a77;
   wire [7:0] _00003a78;
   wire [0:0] _00003a79;
   wire [7:0] _00003a135_00003a_00003areg__0;
   wire [7:0] _00003a135_00003a_00003areg__1;
   wire [0:0] _00003a135_00003a_00003a_00003a120_00003a_00003aabus__r;
   wire [0:0] _00003a135_00003a_00003a_00003a121_00003a_00003aabus__w;
   wire [0:0] _00003a135_00003a_00003a_00003a122_00003a_00003aabus__r;
   wire [0:0] _00003a135_00003a_00003a_00003a123_00003a_00003aabus__w;
   reg [7:0] _00003a136_00003a_00003alv0;
   reg [7:0] _00003a136_00003a_00003alv1;
   reg [7:0] _00003a136_00003a_00003arv0;
   reg [7:0] _00003a136_00003a_00003arv1;
   reg _00003a136_00003a_00003alvok0;
   reg _00003a136_00003a_00003alvok1;
   reg _00003a136_00003a_00003arvok0;
   reg _00003a136_00003a_00003arvok1;
   reg _00003a136_00003a_00003arun;
   wire _00005e_00006060;
   wire _00005e_00006061;

   _____00003aT0_00003a_00003amy__layer_00003aT0_00003a_00003amy__initializer_00003aT0 my__initializer(.clk(_00005e_00006060),.flag(_00005e_00006061));
   assign _00005e_00006060 = clk;

   assign _00005e_00006061 = flag;

   assign _00003a62 = _00003a135_00003a_00003areg__0;

   assign _00003a63 = _00003a135_00003a_00003areg__1;

   assign _00003a77 = _00003a135_00003a_00003areg__0;

   assign _00003a78 = _00003a135_00003a_00003areg__1;

   assign _00003a79 = _00003a135_00003a_00003a_00003a121_00003a_00003aabus__w;

   always @( posedge clk ) begin

      ack <= 32'd0;

      _00003a136_00003a_00003arun <= 32'd0;

      if ((req | _00003a136_00003a_00003arun)) begin
         _00003a136_00003a_00003arun <= 32'd1;
         _00003a136_00003a_00003alv0 <= _00003a2;
         _00003a136_00003a_00003alvok0 <= 32'd1;
         _00003a136_00003a_00003arv0 <= _00003a62;
         _00003a136_00003a_00003arvok0 <= 32'd1;
         if ((_00003a136_00003a_00003alvok0 & _00003a136_00003a_00003arvok0)) begin
            _00003a136_00003a_00003arun <= 32'd0;
            ack <= 32'd1;
            _00003a32 <= (_00003a136_00003a_00003alv0 + _00003a136_00003a_00003arv0);
         end
         _00003a136_00003a_00003alv1 <= _00003a3;
         _00003a136_00003a_00003alvok1 <= 32'd1;
         _00003a136_00003a_00003arv1 <= _00003a63;
         _00003a136_00003a_00003arvok1 <= 32'd1;
         if ((_00003a136_00003a_00003alvok1 & _00003a136_00003a_00003arvok1)) begin
            _00003a136_00003a_00003arun <= 32'd0;
            ack <= 32'd1;
            _00003a33 <= (_00003a136_00003a_00003alv1 + _00003a136_00003a_00003arv1);
         end
      end
      else begin
         _00003a136_00003a_00003alvok0 <= 32'd0;
         _00003a136_00003a_00003arvok0 <= 32'd0;
         _00003a136_00003a_00003alvok1 <= 32'd0;
         _00003a136_00003a_00003arvok1 <= 32'd0;
      end

   end

endmodule